module seven_seg_decoder(SW,LEDR);

		input [1:0]SW;
		output [6:0]LEDR;
		reg u,v,w;

endmodule 